`ifndef UTILS_VH
  `define UTILS_VH

  `define CPU_WSIZE  (8)
  `define CPU_HSIZE  (`CPU_WSIZE>>1)

  // COMMONS:
  `define ZERO       (0)

  // ALU:
  `define ALU_OSIZE  (4)

  `define ALU_AND_OP (0)
  `define ALU_OR_OP  (1)
  `define ALU_ADD_OP (2)
  `define ALU_SUB_OP (6)
  `define ALU_SLT_OP (7)
  `define ALU_LUI_OP (8)
  `define ALU_NOR_OP (12)

  // ALU Control:


`endif // UTILS_VH
